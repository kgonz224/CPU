/*
  Author: Prabakar, FIU-SCIS
   Template for proj4 test bench program
*/

module template_tb; // processor test bench template
  reg [7:0] IMem[4095:0]; // 4096 bytes (1024 words)
  reg [7:0] DMem[8191:0]; // 8192 bytes (1024 double words)
  reg [31:0] instruction; // all instructions are 32-bit wide
  reg [63:0] PC; // PC contains 64-bit byte address

  initial // load instruction memory and data memory
  begin 
	$readmemh("IM_Bytes.txt", IMem);
	$readmemh("DM_Bytes.txt", DMem);
	PC <= 64'b0; // initialize PC
  end 
  
  always //sequential logic of fetch for illustration
  begin
	#1
	// this code block can be performed in any other module
	// concatenate four bytes of IMem into PC
	instruction[7:0] = IMem[PC];
	instruction[15:8] = IMem[PC + 1];
	instruction[23:16] = IMem[PC + 2];
	instruction[31:24] = IMem[PC + 3];
	$display("Opcode value: %11b \n", instruction[31:21]);
	PC = PC + 4; // PC needs to be updated in the processor/datapath module
  end

  // output data memory to a file when HALT instruction is fetched
  always @(instruction) 
  begin
    if (instruction[31:21] == {11{1'b1}})
    begin
	$display("final opcode is detected \n");
	$writememh("DM_Final_Bytes.txt", DMem);
	$finish;
    end
  end
endmodule 
