`include "Execution.v"
`include "CPU_control.v"

module InstructionDecode(InstructionI, AddressI, PCSrc, BranchAddress);

  reg [63:0] Regs [31:0]; // 32 double words
  input [31:0] InstructionI;
  input [63:0] AddressI;
  output PCSrc;
  output [63:0] BranchAddress;
  reg [63:0] Address, Data1, Data2, signExtInstr, AddressO, Data1O, Data2O,
	  signExtInstrO;
  reg [31:0] Instruction, InstructionO;
  reg RegWriteO, BO, BZO, BNZO, MemReadO, MemWriteO, MemtoRegO;
  wire Reg2Loc, RegWrite, B, BZ, BNZ, MemRead, MemWrite, MemtoReg, PCSrc;
  wire [1:0] ALUOp, ALUSrc;
  reg [1:0] ALUOpO, ALUSrcO;

  initial
  begin
	Regs[31] = {64{1'b0}};
	Instruction = {32{1'b0}};
  end

  cpu_control controlUnit(Instruction[31:21], Reg2Loc, B, BZ, BNZ,
	  MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc, RegWrite);

  
  Execution ex(AddressO, InstructionO, signExtInstrO, Data1O, Data2O, ALUSrcO,
	  ALUOpO, BO, BZO, BNZO, MemWriteO, MemReadO, MemtoRegO, RegWriteO,
	  Data2Write, Reg2Write, OldRegWrite, BranchAddress, PCSrc);

always
  begin
	  #1
	  Address = AddressI;
	  Instruction = InstructionI;
	  #2;
  end

always@(Instruction)
  begin
	  $display("IDcode value: %32b %d\n", Instruction[31:0], $time);
	  Data1 <= Regs[Instruction[9:5]];
	  #1
	  if (Reg2Loc == 0)
	          Data2 = Regs[Instruction[20:16]];
	  else
                  Data2[7:0] = Regs[Instruction[4:0]];

	  if(B)
	  begin
		  signExtInstr[25:0] = Instruction[25:0];
		  signExtInstr[63:45] = {38{Instruction[25]}};  
	  end
	  else if(BZ | BNZ)
	  begin		  
		  signExtInstr[18:0] = Instruction[23:5];
		  signExtInstr[63:45] = {45{Instruction[23]}};
	  end
	  else
	  begin
		  signExtInstr[9:0] = Instruction[20:11];
		  signExtInstr[63:10] = {54{Instruction[20]}};
	  end

  end

  always
  begin
	#3
  	AddressO = Address;
        Data1O = Data1;
       	Data2O = Data2;
       	signExtInstrO = signExtInstr;
	ALUSrcO = ALUSrc;
	ALUOpO = ALUOp;
       	RegWriteO = RegWrite;
       	BO = B; 
	BZO = BZ;
	BNZO = BNZ;
       	MemReadO = MemRead;
	MemWriteO = MemWrite;
       	MemtoRegO = MemtoReg;
        InstructionO = InstructionO;
  end

  always @(OldRegWrite)
  begin
	Regs[Reg2Write] = Data2Write;
  end
endmodule

